module wire(output out, input in);
    assign out = in;
endmodule